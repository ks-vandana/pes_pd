* SPICE3 file created from sky130_inv.ext - technology: sky130A

.option scale=10000u

.subckt sky130_inv A Y VPWR VGND
M1000 Y A VPWR VPWR pshort w=37 l=23
+  ad=1443 pd=152 as=1517 ps=156
M1001 Y A VGND VGND nshort w=35 l=23
+  ad=1435 pd=152 as=1365 ps=148
C0 A VPWR 0.07fF
C1 VPWR Y 0.11fF
C2 A Y 0.05fF
C3 Y VGND 0.24fF
C4 VPWR VGND 0.59fF
.ends
